library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity bit_feeder is
    Port (
        clk        : in  std_logic;
        reset      : in  std_logic;
        bit_out    : out std_logic;
        strobe_out : out std_logic
    );
end entity;

architecture bit_feeder_arch of bit_feeder is

    constant ROM_SIZE : integer := 2048;

    type rom_type is array (0 to ROM_SIZE - 1) of std_logic_vector(1 downto 0);
    constant rom : rom_type := (
		0 => "00", 1 => "00", 2 => "00", 3 => "00", 4 => "00", 5 => "00", 6 => "00", 7 => "00", 8 => "00", 9 => "00", 10 => "00", 11 => "00", 12 => "00", 13 => "00", 14 => "00", 15 => "00", 16 => "00", 17 => "00", 18 => "00", 19 => "00", 20 => "00", 21 => "00", 22 => "00", 23 => "00", 24 => "00", 25 => "00", 26 => "00", 27 => "00", 28 => "00", 29 => "00", 30 => "00", 31 => "00", 32 => "00", 33 => "00", 34 => "00", 35 => "00", 36 => "00", 37 => "00", 38 => "00", 39 => "00", 40 => "00", 41 => "00", 42 => "00", 43 => "00", 44 => "00", 45 => "00", 46 => "00", 47 => "00", 48 => "00", 49 => "00", 50 => "00", 51 => "00", 52 => "00", 53 => "00", 54 => "00", 55 => "00", 56 => "00", 57 => "00", 58 => "00", 59 => "00", 60 => "00", 61 => "00", 62 => "00", 63 => "00", 64 => "00", 65 => "00", 66 => "00", 67 => "00", 68 => "00", 69 => "00", 70 => "00", 71 => "00", 72 => "00", 73 => "00", 74 => "00", 75 => "00", 76 => "00", 77 => "00", 78 => "00", 79 => "00", 80 => "00", 81 => "00", 82 => "00", 83 => "00", 84 => "00", 85 => "00", 86 => "00", 87 => "00", 88 => "00", 89 => "00", 90 => "00", 91 => "00", 92 => "00", 93 => "00", 94 => "00", 95 => "00", 96 => "00", 97 => "00", 98 => "00", 99 => "00", 100 => "00", 101 => "00", 102 => "00", 103 => "00", 104 => "00", 105 => "00", 106 => "00", 107 => "00", 108 => "00", 109 => "00", 110 => "00", 111 => "00", 112 => "00", 113 => "00", 114 => "00", 115 => "00", 116 => "00", 117 => "00", 118 => "00", 119 => "00", 120 => "00", 121 => "00", 122 => "00", 123 => "00", 124 => "00", 125 => "00", 126 => "00", 127 => "00", 128 => "00", 129 => "00", 130 => "00", 131 => "00", 132 => "00", 133 => "00", 134 => "00", 135 => "00", 136 => "00", 137 => "00", 138 => "00", 139 => "00", 140 => "00", 141 => "00", 142 => "00", 143 => "00", 144 => "00", 145 => "00", 146 => "00", 147 => "00", 148 => "00", 149 => "00", 150 => "00", 151 => "00", 152 => "00", 153 => "00", 154 => "00", 155 => "00", 156 => "00", 157 => "00", 158 => "00", 159 => "00", 160 => "00", 161 => "00", 162 => "00", 163 => "00", 164 => "00", 165 => "00", 166 => "00", 167 => "00", 168 => "00", 169 => "00", 170 => "00", 171 => "00", 172 => "00", 173 => "00", 174 => "00", 175 => "00", 176 => "00", 177 => "00", 178 => "00", 179 => "00", 180 => "00", 181 => "00", 182 => "00", 183 => "00", 184 => "00", 185 => "00", 186 => "00", 187 => "00", 188 => "00", 189 => "00", 190 => "00", 191 => "00", 192 => "00", 193 => "00", 194 => "00", 195 => "00", 196 => "00", 197 => "00", 198 => "00", 199 => "00", 200 => "00", 201 => "00", 202 => "00", 203 => "00", 204 => "00", 205 => "00", 206 => "00", 207 => "00", 208 => "00", 209 => "00", 210 => "00", 211 => "00", 212 => "00", 213 => "00", 214 => "00", 215 => "00", 216 => "00", 217 => "00", 218 => "00", 219 => "00", 220 => "00", 221 => "00", 222 => "00", 223 => "00", 224 => "00", 225 => "00", 226 => "00", 227 => "00", 228 => "00", 229 => "00", 230 => "00", 231 => "00", 232 => "00", 233 => "00", 234 => "00", 235 => "00", 236 => "00", 237 => "00", 238 => "00", 239 => "00", 240 => "00", 241 => "00", 242 => "00", 243 => "00", 244 => "00", 245 => "00", 246 => "00", 247 => "00", 248 => "00", 249 => "00", 250 => "00", 251 => "00", 252 => "00", 253 => "00", 254 => "00", 255 => "00", 256 => "00", 257 => "00", 258 => "00", 259 => "00", 260 => "00", 261 => "00", 262 => "00", 263 => "00", 264 => "00", 265 => "00", 266 => "00", 267 => "00", 268 => "00", 269 => "00", 270 => "00", 271 => "00", 272 => "00", 273 => "00", 274 => "00", 275 => "00", 276 => "00", 277 => "00", 278 => "00", 279 => "00", 280 => "00", 281 => "00", 282 => "00", 283 => "00", 284 => "00", 285 => "00", 286 => "00", 287 => "00", 288 => "00", 289 => "00", 290 => "00", 291 => "00", 292 => "00", 293 => "00", 294 => "00", 295 => "00", 296 => "00", 297 => "00", 298 => "00", 299 => "00", 300 => "00", 301 => "00", 302 => "00", 303 => "00", 304 => "00", 305 => "00", 306 => "00", 307 => "00", 308 => "00", 309 => "00", 310 => "00", 311 => "00", 312 => "00", 313 => "00", 314 => "00", 315 => "00", 316 => "00", 317 => "00", 318 => "00", 319 => "00", 320 => "00", 321 => "00", 322 => "00", 323 => "00", 324 => "00", 325 => "00", 326 => "00", 327 => "00", 328 => "00", 329 => "00", 330 => "00", 331 => "00", 332 => "00", 333 => "00", 334 => "00", 335 => "00", 336 => "00", 337 => "00", 338 => "00", 339 => "00", 340 => "00", 341 => "00", 342 => "00", 343 => "00", 344 => "00", 345 => "00", 346 => "00", 347 => "00", 348 => "00", 349 => "00", 350 => "00", 351 => "00", 352 => "00", 353 => "00", 354 => "00", 355 => "00", 356 => "00", 357 => "00", 358 => "00", 359 => "00", 360 => "00", 361 => "00", 362 => "00", 363 => "00", 364 => "00", 365 => "00", 366 => "00", 367 => "00", 368 => "00", 369 => "00", 370 => "00", 371 => "00", 372 => "00", 373 => "00", 374 => "00", 375 => "00", 376 => "00", 377 => "00", 378 => "00", 379 => "00", 380 => "00", 381 => "00", 382 => "00", 383 => "00", 384 => "00", 385 => "00", 386 => "00", 387 => "00", 388 => "00", 389 => "00", 390 => "00", 391 => "00", 392 => "00", 393 => "00", 394 => "00", 395 => "00", 396 => "00", 397 => "00", 398 => "00", 399 => "00", 400 => "00", 401 => "00", 402 => "00", 403 => "00", 404 => "00", 405 => "00", 406 => "00", 407 => "00", 408 => "00", 409 => "00", 410 => "00", 411 => "00", 412 => "00", 413 => "00", 414 => "00", 415 => "00", 416 => "00", 417 => "00", 418 => "00", 419 => "00", 420 => "00", 421 => "00", 422 => "00", 423 => "00", 424 => "00", 425 => "00", 426 => "00", 427 => "00", 428 => "00", 429 => "00", 430 => "00", 431 => "00", 432 => "00", 433 => "00", 434 => "00", 435 => "00", 436 => "00", 437 => "00", 438 => "00", 439 => "00", 440 => "00", 441 => "00", 442 => "00", 443 => "00", 444 => "00", 445 => "00", 446 => "00", 447 => "00", 448 => "00", 449 => "00", 450 => "00", 451 => "00", 452 => "00", 453 => "00", 454 => "00", 455 => "00", 456 => "00", 457 => "00", 458 => "00", 459 => "00", 460 => "00", 461 => "00", 462 => "00", 463 => "00", 464 => "00", 465 => "00", 466 => "00", 467 => "00", 468 => "00", 469 => "00", 470 => "00", 471 => "00", 472 => "00", 473 => "00", 474 => "00", 475 => "00", 476 => "00", 477 => "00", 478 => "00", 479 => "00", 480 => "00", 481 => "00", 482 => "00", 483 => "00", 484 => "00", 485 => "00", 486 => "00", 487 => "00", 488 => "00", 489 => "00", 490 => "00", 491 => "00", 492 => "00", 493 => "00", 494 => "00", 495 => "00", 496 => "00", 497 => "00", 498 => "00", 499 => "00", 500 => "00", 501 => "00", 502 => "00", 503 => "00", 504 => "00", 505 => "00", 506 => "00", 507 => "00", 508 => "00", 509 => "00", 510 => "00", 511 => "00", 512 => "00", 513 => "00", 514 => "00", 515 => "00", 516 => "00", 517 => "00", 518 => "00", 519 => "00", 520 => "00", 521 => "00", 522 => "00", 523 => "00", 524 => "00", 525 => "00", 526 => "00", 527 => "00", 528 => "00", 529 => "00", 530 => "00", 531 => "00", 532 => "00", 533 => "00", 534 => "00", 535 => "00", 536 => "00", 537 => "00", 538 => "00", 539 => "00", 540 => "00", 541 => "00", 542 => "00", 543 => "00", 544 => "00", 545 => "00", 546 => "00", 547 => "00", 548 => "00", 549 => "00", 550 => "00", 551 => "00", 552 => "00", 553 => "00", 554 => "00", 555 => "00", 556 => "00", 557 => "00", 558 => "00", 559 => "00", 560 => "00", 561 => "00", 562 => "00", 563 => "00", 564 => "00", 565 => "00", 566 => "00", 567 => "00", 568 => "00", 569 => "00", 570 => "00", 571 => "00", 572 => "00", 573 => "00", 574 => "00", 575 => "00", 576 => "00", 577 => "00", 578 => "00", 579 => "00", 580 => "00", 581 => "00", 582 => "00", 583 => "00", 584 => "00", 585 => "00", 586 => "00", 587 => "00", 588 => "00", 589 => "00", 590 => "00", 591 => "00", 592 => "00", 593 => "00", 594 => "00", 595 => "00", 596 => "00", 597 => "00", 598 => "00", 599 => "00", 600 => "00", 601 => "00", 602 => "00", 603 => "00", 604 => "00", 605 => "00", 606 => "00", 607 => "00", 608 => "00", 609 => "00", 610 => "00", 611 => "00", 612 => "00", 613 => "00", 614 => "00", 615 => "00", 616 => "00", 617 => "00", 618 => "00", 619 => "00", 620 => "00", 621 => "00", 622 => "00", 623 => "00", 624 => "00", 625 => "00", 626 => "00", 627 => "00", 628 => "00", 629 => "00", 630 => "00", 631 => "00", 632 => "00", 633 => "00", 634 => "00", 635 => "00", 636 => "00", 637 => "00", 638 => "00", 639 => "00", 640 => "00", 641 => "00", 642 => "00", 643 => "00", 644 => "00", 645 => "00", 646 => "00", 647 => "00", 648 => "00", 649 => "00", 650 => "00", 651 => "00", 652 => "00", 653 => "00", 654 => "00", 655 => "00", 656 => "00", 657 => "00", 658 => "00", 659 => "00", 660 => "00", 661 => "00", 662 => "00", 663 => "00", 664 => "00", 665 => "00", 666 => "00", 667 => "00", 668 => "00", 669 => "00", 670 => "00", 671 => "00", 672 => "00", 673 => "00", 674 => "00", 675 => "00", 676 => "00", 677 => "00", 678 => "00", 679 => "00", 680 => "00", 681 => "00", 682 => "00", 683 => "00", 684 => "00", 685 => "00", 686 => "00", 687 => "00", 688 => "00", 689 => "00", 690 => "00", 691 => "00", 692 => "00", 693 => "00", 694 => "00", 695 => "00", 696 => "00", 697 => "00", 698 => "00", 699 => "00", 700 => "00", 701 => "00", 702 => "00", 703 => "00", 704 => "00", 705 => "00", 706 => "00", 707 => "00", 708 => "00", 709 => "00", 710 => "00", 711 => "00", 712 => "00", 713 => "00", 714 => "00", 715 => "00", 716 => "00", 717 => "00", 718 => "00", 719 => "00", 720 => "00", 721 => "00", 722 => "00", 723 => "00", 724 => "00", 725 => "00", 726 => "00", 727 => "00", 728 => "00", 729 => "00", 730 => "00", 731 => "00", 732 => "00", 733 => "00", 734 => "00", 735 => "00", 736 => "00", 737 => "00", 738 => "00", 739 => "00", 740 => "00", 741 => "00", 742 => "00", 743 => "00", 744 => "00", 745 => "00", 746 => "00", 747 => "00", 748 => "00", 749 => "00", 750 => "00", 751 => "00", 752 => "00", 753 => "00", 754 => "00", 755 => "00", 756 => "00", 757 => "00", 758 => "00", 759 => "00", 760 => "00", 761 => "00", 762 => "00", 763 => "00", 764 => "00", 765 => "00", 766 => "00", 767 => "00", 768 => "00", 769 => "00", 770 => "00", 771 => "00", 772 => "00", 773 => "00", 774 => "00", 775 => "00", 776 => "00", 777 => "00", 778 => "00", 779 => "00", 780 => "00", 781 => "00", 782 => "00", 783 => "00", 784 => "00", 785 => "00", 786 => "00", 787 => "00", 788 => "00", 789 => "00", 790 => "00", 791 => "00", 792 => "00", 793 => "00", 794 => "00", 795 => "00", 796 => "00", 797 => "00", 798 => "00", 799 => "00", 800 => "00", 801 => "00", 802 => "00", 803 => "00", 804 => "00", 805 => "00", 806 => "00", 807 => "00", 808 => "00", 809 => "00", 810 => "00", 811 => "00", 812 => "00", 813 => "00", 814 => "00", 815 => "00", 816 => "00", 817 => "00", 818 => "00", 819 => "00", 820 => "00", 821 => "00", 822 => "00", 823 => "00", 824 => "00", 825 => "00", 826 => "00", 827 => "00", 828 => "00", 829 => "00", 830 => "00", 831 => "00", 832 => "00", 833 => "00", 834 => "00", 835 => "00", 836 => "00", 837 => "00", 838 => "00", 839 => "00", 840 => "00", 841 => "00", 842 => "00", 843 => "00", 844 => "00", 845 => "00", 846 => "00", 847 => "00", 848 => "00", 849 => "00", 850 => "00", 851 => "00", 852 => "00", 853 => "00", 854 => "00", 855 => "00", 856 => "00", 857 => "00", 858 => "00", 859 => "00", 860 => "00", 861 => "00", 862 => "00", 863 => "00", 864 => "00", 865 => "00", 866 => "00", 867 => "00", 868 => "00", 869 => "00", 870 => "00", 871 => "00", 872 => "00", 873 => "00", 874 => "00", 875 => "00", 876 => "00", 877 => "00", 878 => "00", 879 => "00", 880 => "00", 881 => "00", 882 => "00", 883 => "00", 884 => "00", 885 => "00", 886 => "00", 887 => "00", 888 => "00", 889 => "00", 890 => "00", 891 => "00", 892 => "00", 893 => "00", 894 => "00", 895 => "00", 896 => "00", 897 => "00", 898 => "00", 899 => "00", 900 => "00", 901 => "00", 902 => "00", 903 => "00", 904 => "00", 905 => "00", 906 => "00", 907 => "00", 908 => "00", 909 => "00", 910 => "00", 911 => "00", 912 => "00", 913 => "00", 914 => "00", 915 => "00", 916 => "00", 917 => "00", 918 => "00", 919 => "00", 920 => "00", 921 => "00", 922 => "00", 923 => "00", 924 => "00", 925 => "00", 926 => "00", 927 => "00", 928 => "00", 929 => "00", 930 => "00", 931 => "00", 932 => "00", 933 => "00", 934 => "00", 935 => "00", 936 => "00", 937 => "00", 938 => "00", 939 => "00", 940 => "00", 941 => "00", 942 => "00", 943 => "00", 944 => "00", 945 => "00", 946 => "00", 947 => "00", 948 => "00", 949 => "00", 950 => "00", 951 => "00", 952 => "00", 953 => "00", 954 => "00", 955 => "00", 956 => "00", 957 => "00", 958 => "00", 959 => "00", 960 => "01", 961 => "11", 962 => "10", 963 => "11", 964 => "01", 965 => "11", 966 => "01", 967 => "00", 968 => "10", 969 => "11", 970 => "10", 971 => "11", 972 => "01", 973 => "11", 974 => "01", 975 => "00", 976 => "10", 977 => "11", 978 => "10", 979 => "11", 980 => "01", 981 => "11", 982 => "01", 983 => "00", 984 => "10", 985 => "11", 986 => "10", 987 => "11", 988 => "01", 989 => "11", 990 => "01", 991 => "00", 992 => "10", 993 => "11", 994 => "10", 995 => "11", 996 => "01", 997 => "11", 998 => "01", 999 => "00", 1000 => "10", 1001 => "11", 1002 => "10", 1003 => "11", 1004 => "01", 1005 => "11", 1006 => "01", 1007 => "00", 1008 => "10", 1009 => "11", 1010 => "10", 1011 => "11", 1012 => "01", 1013 => "11", 1014 => "01", 1015 => "00", 1016 => "10", 1017 => "11", 1018 => "10", 1019 => "11", 1020 => "01", 1021 => "11", 1022 => "01", 1023 => "00", 1024 => "10", 1025 => "11", 1026 => "10", 1027 => "11", 1028 => "01", 1029 => "11", 1030 => "01", 1031 => "00", 1032 => "10", 1033 => "11", 1034 => "10", 1035 => "11", 1036 => "01", 1037 => "11", 1038 => "01", 1039 => "00", 1040 => "10", 1041 => "11", 1042 => "10", 1043 => "11", 1044 => "01", 1045 => "11", 1046 => "01", 1047 => "00", 1048 => "10", 1049 => "11", 1050 => "01", 1051 => "00", 1052 => "10", 1053 => "00", 1054 => "01", 1055 => "11", 1056 => "01", 1057 => "00", 1058 => "10", 1059 => "00", 1060 => "01", 1061 => "00", 1062 => "10", 1063 => "00", 1064 => "01", 1065 => "11", 1066 => "10", 1067 => "00", 1068 => "01", 1069 => "11", 1070 => "01", 1071 => "11", 1072 => "10", 1073 => "00", 1074 => "01", 1075 => "11", 1076 => "10", 1077 => "00", 1078 => "10", 1079 => "11", 1080 => "01", 1081 => "00", 1082 => "10", 1083 => "00", 1084 => "01", 1085 => "11", 1086 => "10", 1087 => "00", 1088 => "10", 1089 => "11", 1090 => "01", 1091 => "00", 1092 => "10", 1093 => "00", 1094 => "01", 1095 => "11", 1096 => "10", 1097 => "00", 1098 => "10", 1099 => "11", 1100 => "10", 1101 => "11", 1102 => "10", 1103 => "00", 1104 => "01", 1105 => "00", 1106 => "10", 1107 => "00", 1108 => "01", 1109 => "00", 1110 => "01", 1111 => "00", 1112 => "01", 1113 => "00", 1114 => "01", 1115 => "11", 1116 => "01", 1117 => "11", 1118 => "01", 1119 => "11", 1120 => "10", 1121 => "11", 1122 => "01", 1123 => "00", 1124 => "01", 1125 => "11", 1126 => "10", 1127 => "00", 1128 => "10", 1129 => "11", 1130 => "10", 1131 => "11", 1132 => "10", 1133 => "00", 1134 => "01", 1135 => "11", 1136 => "10", 1137 => "11", 1138 => "01", 1139 => "00", 1140 => "10", 1141 => "00", 1142 => "10", 1143 => "00", 1144 => "01", 1145 => "11", 1146 => "10", 1147 => "00", 1148 => "01", 1149 => "11", 1150 => "01", 1151 => "00", 1152 => "10", 1153 => "11", 1154 => "01", 1155 => "11", others => "00");
    signal address			: integer range 0 to ROM_SIZE - 1 := 0;

begin
    process(clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                address     		<= 0;
            else
                bit_out		<= rom(address)(1);
					 strobe_out	<= rom(address)(0);
                address		<= address + 1;
            end if;
        end if;
    end process;
end architecture;